module exercise24
(
	input logic clk, reset,
	input logic a, b,
	output logic y
);
	logic [1:0] state, nextstate;
	parameter S0 = 2'b00;
	parameter S1 = 2'b01;
	parameter S2 = 2'b10;
	parameter S3 = 2'b11;
	always_ff @(posedge clk, posedge reset)
		if (reset) state <= S0;
		else	   state <= nextstate;
		always_comb
			case(state)
				S0: if (a ^ b) nextstate = S1;
					else	   nextstate = S0;
				S1: if (a & b) nextstate = S2;
					else 	   nextstate = S0;
				S2: if (a | b) nextstate = S3;
					else	   nextstate = S0;
				S3: if (a | b) nextstate = S3;
					else	   nextstate = S0;
			endcase
		assign y = (state == S1) | (state == S2);
endmodule
