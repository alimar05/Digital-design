module testbench1();
	logic a, b, c, y;
	// instantiate device under test
	example dut(a, b, c, y);
	// apply unputs one at a time
	initial begin
		a = 0; b = 0; c = 0; #10;
		c = 1; 		     #10;
		b = 1; c = 0;        #10;
		c = 1; 		     #10;
		a = 1; b = 0; c = 0; #10;
		c = 1; 		     #10;
		b = 1; c = 0; 	     #10;
		c = 1; 		     #10;
	 end
endmodule
