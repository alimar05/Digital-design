module exercise19
(
	input logic [3:0] a,
	output logic p, d
);
	always_comb
		case(a)
			0: {p, d} = 2'b00;
			1: {p, d} = 2'b00;
			2: {p, d} = 2'b10;
			3: {p, d} = 2'b11;
			4: {p, d} = 2'b00;
			5: {p, d} = 2'b10;
			6: {p, d} = 2'b01;
			7: {p, d} = 2'b10;
			8: {p, d} = 2'b00;
			9: {p, d} = 2'b01;
		   10: {p, d} = 2'b00;
		   11: {p, d} = 2'b10;
	       12: {p, d} = 2'b01;
		   13: {p, d} = 2'b10;
		   14: {p, d} = 2'b00;
		   15: {p, d} = 2'b01;
		endcase
endmodule
